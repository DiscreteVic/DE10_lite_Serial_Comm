// unsaved.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module unsaved (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	unsaved_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),        //          clk.clk
		.clk_reset_reset      (~reset_reset_n), //    clk_reset.reset
		.master_address       (),               //       master.address
		.master_readdata      (),               //             .readdata
		.master_read          (),               //             .read
		.master_write         (),               //             .write
		.master_writedata     (),               //             .writedata
		.master_waitrequest   (),               //             .waitrequest
		.master_readdatavalid (),               //             .readdatavalid
		.master_byteenable    (),               //             .byteenable
		.master_reset_reset   ()                // master_reset.reset
	);

endmodule
